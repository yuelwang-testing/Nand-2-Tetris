module Not(
  input in,
  output out
);
  nand gate1(out, in, in);
endmodule
